assign o_d_conn_<i_pre>C<i_post>[<i_dim>] = uart_rx_data[<bit_post> : <bit_pre>];
    <rx-flag>