    assign i_d_ensemble_<i_post>[<current_i>] = o_d_conn_<i_pre>C<i_post>;
    assign i_d_valids_<i_post>[<current_i>] = o_d_valid_conn_<i_pre>C<i_post>;