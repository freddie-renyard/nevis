    /**************** CONNECTION 0C<i_pre>+N *************/
    wire [OUTPUT_DIMS_<i_pre>C<i_post>-1:0][N_OUTPUT_<i_pre>C<i_post>-1:0]    o_output_val;
    wire [OUTPUT_DIMS_<i_pre>C<i_post>-1:0]                      o_output_valid;

