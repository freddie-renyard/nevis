    assign o_d_valid_conn_<i_pre>C<i_post> = o_scheduler;
