    /**************** CONNECTION <i_pre>C<i_post> WIRES *************/
    wire [OUTPUT_DIMS_<i_pre>C<i_post>-1:0][N_OUTPUT_<i_pre>C<i_post>-1:0] o_d_conn_<i_pre>C<i_post>;
    wire [OUTPUT_DIMS_<i_pre>C<i_post>-1:0] o_d_valid_conn_<i_pre>C<i_post>;

