    assign i_d_ensemble_<i_pre>[<current_i>] = o_d_conn_<i_pre>C<i_post>
