    assign i_d_valids_<i_post>[<current_i>] = o_d_valid_conn_<i_pre>C<i_post>;
    