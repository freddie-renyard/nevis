    assign i_d_ensemble_<i_post>[<current_dim>][<current_i>] = o_d_conn_<i_pre>C<i_post>[<current_dim>];
