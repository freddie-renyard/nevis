assign uart_tx_data[<bit_post> : <bit_pre>] = o_d_conn_<i_pre>C<i_post>[<i_dim>];
    <tx-flag>