    assign i_d_valids_<i>[<input_index>] = o_d_valid_conn_<i_pre>C<i>;

