// Population A Params
parameter N_NEURON_A = 50,
N_X_A = 8,
RADIX_X_A = 7,
N_G_MAN_A = 7,
N_G_EXP_A = 4,
N_B_MAN_A = 7,
N_B_EXP_A = 4,
N_DV_POST_A = 10;

// Population A Synaptic Params
parameter N_WEIGHT_A = 16,
SCALE_W_A = 5,
N_WEIGHT_EXP_A = 5,
N_ACTIV_EXTRA_A = 6,
PSTC_SHIFT_A = 7;

// Population B Params
parameter N_NEURON_B = 40,
N_X_B = 23,
RADIX_X_B = 21,
N_G_MAN_B = 7,
N_G_EXP_B = 4,
N_B_MAN_B = 7,
N_B_EXP_B = 4,
N_DV_POST_B = 10;

// Population B Synaptic Params
parameter N_WEIGHT_B = 16,
SCALE_W_B = 6,
N_WEIGHT_EXP_B = 5,
N_ACTIV_EXTRA_B = 8,
PSTC_SHIFT_B = 7;

// Global Synaptic Params
parameter N_R = 2,
REF_VALUE = 1,
T_RC_SHIFT = 4;
